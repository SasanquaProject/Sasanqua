module decode_1
    (
        /* ----- 制御 ----- */
        input wire          CLK,
        input wire          RST
    );

endmodule
