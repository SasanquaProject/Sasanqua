module mmu
    (
    );

endmodule
