module decode_2
    (
        /* ----- 制御 ----- */
        input wire          CLK,
        input wire          RST
    );

endmodule
