module core
    (
        /* ----- 制御 ----- */
        input wire          CLK,
        input wire          RST,

        /* ----- メモリアクセス信号 ----- */
        // 命令
        output reg          INST_RDEN,
        output reg  [31:0]  INST_RADDR,
        input wire          INST_RVALID,
        input wire  [31:0]  INST_RDATA,

        // データ
        // input wire          DATA_WREN,
        // input wire [31:0]   DATA_WRADDR,
        // input wire [31:0]   DATA_WRDATA,
        output wire         DATA_RDEN,
        output wire [31:0]  DATA_RADDR,
        input wire          DATA_RVALID,
        input wire  [31:0]  DATA_RDATA,

        // ハザード
        input wire          MEM_WAIT
    );

    assign DATA_RDEN    = 1'b0;
    assign DATA_RADDR   = 32'b0;

    /* ----- 1. 命令フェッチ ----- */
    wire        inst_valid;
    wire [31:0] inst_addr, inst_data;

    assign inst_valid   = INST_RVALID;
    assign inst_addr    = INST_RADDR;
    assign inst_data    = INST_RDATA;

    always @ (posedge CLK) begin
        if (RST) begin
            INST_RDEN <= 1'b0;
            INST_RADDR <= 32'hffff_fffc;
        end
        else if (!MEM_WAIT) begin
            INST_RDEN <= 1'b1;
            INST_RADDR <= INST_RADDR + 32'd4;
        end
    end

    /* ----- 2. 命令デコード1 ----- */
    wire        decode_1st_valid;
    wire [31:0] decode_1st_pc, decode_1st_imm_i, decode_1st_imm_s, decode_1st_imm_b, decode_1st_imm_u, decode_1st_imm_j;
    wire [6:0]  decode_1st_opcode, decode_1st_funct7;
    wire [4:0]  decode_1st_rd, decode_1st_rs1, decode_1st_rs2;
    wire [2:0]  decode_1st_funct3;

    decode_1st decode_1st (
        // 制御
        .CLK            (CLK),
        .RST            (RST),

        // フェッチ部との接続
        .INST_VALID     (inst_valid),
        .INST_PC        (inst_addr),
        .INST_DATA      (inst_data),

        // デコード部2との接続
        .DECODE_1ST_VALID  (decode_1st_valid),
        .DECODE_1ST_PC     (decode_1st_pc),
        .DECODE_1ST_OPCODE (decode_1st_opcode),
        .DECODE_1ST_RD     (decode_1st_rd),
        .DECODE_1ST_RS1    (decode_1st_rs1),
        .DECODE_1ST_RS2    (decode_1st_rs2),
        .DECODE_1ST_FUNCT3 (decode_1st_funct3),
        .DECODE_1ST_FUNCT7 (decode_1st_funct7),
        .DECODE_1ST_IMM_I  (decode_1st_imm_i),
        .DECODE_1ST_IMM_S  (decode_1st_imm_s),
        .DECODE_1ST_IMM_B  (decode_1st_imm_b),
        .DECODE_1ST_IMM_U  (decode_1st_imm_u),
        .DECODE_1ST_IMM_J  (decode_1st_imm_j)
    );

    /* ----- 3. 命令デコード2 ----- */
    wire        decode_2nd_valid;
    wire [31:0] decode_2nd_pc, decode_2nd_imm;
    wire [6:0]  decode_2nd_opcode, decode_2nd_funct7;
    wire [4:0]  decode_2nd_rd, decode_2nd_rs1, decode_2nd_rs2;
    wire [2:0]  decode_2nd_funct3;

    decode_2nd decode_2nd (
        // 制御
        .CLK            (CLK),
        .RST            (RST),

        // デコード部1との接続
        .DECODE_1ST_VALID  (decode_1st_valid),
        .DECODE_1ST_PC     (decode_1st_pc),
        .DECODE_1ST_OPCODE (decode_1st_opcode),
        .DECODE_1ST_RD     (decode_1st_rd),
        .DECODE_1ST_RS1    (decode_1st_rs1),
        .DECODE_1ST_RS2    (decode_1st_rs2),
        .DECODE_1ST_FUNCT3 (decode_1st_funct3),
        .DECODE_1ST_FUNCT7 (decode_1st_funct7),
        .DECODE_1ST_IMM_I  (decode_1st_imm_i),
        .DECODE_1ST_IMM_S  (decode_1st_imm_s),
        .DECODE_1ST_IMM_B  (decode_1st_imm_b),
        .DECODE_1ST_IMM_U  (decode_1st_imm_u),
        .DECODE_1ST_IMM_J  (decode_1st_imm_j),

        .DECODE_2ND_VALID  (decode_2nd_valid),
        .DECODE_2ND_PC     (decode_2nd_pc),
        .DECODE_2ND_OPCODE (decode_2nd_opcode),
        .DECODE_2ND_RD     (decode_2nd_rd),
        .DECODE_2ND_RS1    (decode_2nd_rs1),
        .DECODE_2ND_RS2    (decode_2nd_rs2),
        .DECODE_2ND_FUNCT3 (decode_2nd_funct3),
        .DECODE_2ND_FUNCT7 (decode_2nd_funct7),
        .DECODE_2ND_IMM    (decode_2nd_imm)
    );

    // /* ----- 3-2. レジスタアクセス ----- */
    // wire [31:0] reg_rs1_v, reg_rs2_v;

    // register register (
    //     // 制御
    //     .CLK        (CLK),
    //     .RST        (RST),

    //     // レジスタアクセス(rv32i)
    //     .REG_IR_A   (decode1_rs1),
    //     .REG_IR_B   (decode1_rs2),
    //     .REG_IR_AV  (reg_rs1_v),
    //     .REG_IR_BV  (reg_rs2_v)
    // );

    /* ----- 4. 実行 ----- */
    exec exec (
        // 制御
        .CLK    (CLK),
        .RST    (RST)
    );

    /* ----- 5. メモリアクセス ----- */


endmodule
