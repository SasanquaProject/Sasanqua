module clint
    (
    );

endmodule
